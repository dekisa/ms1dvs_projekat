-- processor_system.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity processor_system is
	port (
		clk_clk       : in    std_logic                     := '0';             --       clk.clk
		reset_reset_n : in    std_logic                     := '0';             --     reset.reset_n
		sdram_addr    : out   std_logic_vector(12 downto 0);                    --     sdram.addr
		sdram_ba      : out   std_logic_vector(1 downto 0);                     --          .ba
		sdram_cas_n   : out   std_logic;                                        --          .cas_n
		sdram_cke     : out   std_logic;                                        --          .cke
		sdram_cs_n    : out   std_logic;                                        --          .cs_n
		sdram_dq      : inout std_logic_vector(15 downto 0) := (others => '0'); --          .dq
		sdram_dqm     : out   std_logic_vector(1 downto 0);                     --          .dqm
		sdram_ras_n   : out   std_logic;                                        --          .ras_n
		sdram_we_n    : out   std_logic;                                        --          .we_n
		sdram_clk_clk : out   std_logic                                         -- sdram_clk.clk
	);
end entity processor_system;

architecture rtl of processor_system is
	component acc_linear_function is
		port (
			reset                  : in  std_logic                     := 'X';             -- reset
			avs_params_address     : in  std_logic                     := 'X';             -- address
			avs_params_read        : in  std_logic                     := 'X';             -- read
			avs_params_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avs_params_write       : in  std_logic                     := 'X';             -- write
			avs_params_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_params_waitrequest : out std_logic;                                        -- waitrequest
			clk                    : in  std_logic                     := 'X';             -- clk
			asi_in_data            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			asi_in_ready           : out std_logic;                                        -- ready
			asi_in_valid           : in  std_logic                     := 'X';             -- valid
			asi_in_eop             : in  std_logic                     := 'X';             -- endofpacket
			asi_in_sop             : in  std_logic                     := 'X';             -- startofpacket
			aso_out_data           : out std_logic_vector(31 downto 0);                    -- data
			aso_out_ready          : in  std_logic                     := 'X';             -- ready
			aso_out_valid          : out std_logic;                                        -- valid
			aso_out_empty          : out std_logic;                                        -- empty
			aso_out_eop            : out std_logic;                                        -- endofpacket
			aso_out_sop            : out std_logic                                         -- startofpacket
		);
	end component acc_linear_function;

	component processor_system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component processor_system_jtag_uart_0;

	component processor_system_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component processor_system_nios2_gen2_0;

	component processor_system_performance_counter_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component processor_system_performance_counter_0;

	component processor_system_pll is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component processor_system_pll;

	component processor_system_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component processor_system_sdram;

	component processor_system_sgdma_mm2s is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			m_read_readdata               : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			m_read_readdatavalid          : in  std_logic                     := 'X';             -- readdatavalid
			m_read_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			m_read_address                : out std_logic_vector(31 downto 0);                    -- address
			m_read_read                   : out std_logic;                                        -- read
			out_data                      : out std_logic_vector(7 downto 0);                     -- data
			out_valid                     : out std_logic;                                        -- valid
			out_ready                     : in  std_logic                     := 'X';             -- ready
			out_endofpacket               : out std_logic;                                        -- endofpacket
			out_startofpacket             : out std_logic                                         -- startofpacket
		);
	end component processor_system_sgdma_mm2s;

	component processor_system_sgdma_s2mm is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			in_startofpacket              : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket                : in  std_logic                     := 'X';             -- endofpacket
			in_data                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_valid                      : in  std_logic                     := 'X';             -- valid
			in_ready                      : out std_logic;                                        -- ready
			in_empty                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			m_write_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			m_write_address               : out std_logic_vector(31 downto 0);                    -- address
			m_write_write                 : out std_logic;                                        -- write
			m_write_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			m_write_byteenable            : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component processor_system_sgdma_s2mm;

	component processor_system_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                         : in  std_logic                     := 'X';             -- clk
			pll_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset        : in  std_logic                     := 'X';             -- reset
			pll_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                      : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                  : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                         : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                     : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                        : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                  : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address               : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                  : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			sgdma_mm2s_descriptor_read_address                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_mm2s_descriptor_read_waitrequest                : out std_logic;                                        -- waitrequest
			sgdma_mm2s_descriptor_read_read                       : in  std_logic                     := 'X';             -- read
			sgdma_mm2s_descriptor_read_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			sgdma_mm2s_descriptor_read_readdatavalid              : out std_logic;                                        -- readdatavalid
			sgdma_mm2s_descriptor_write_address                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_mm2s_descriptor_write_waitrequest               : out std_logic;                                        -- waitrequest
			sgdma_mm2s_descriptor_write_write                     : in  std_logic                     := 'X';             -- write
			sgdma_mm2s_descriptor_write_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sgdma_mm2s_m_read_address                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_mm2s_m_read_waitrequest                         : out std_logic;                                        -- waitrequest
			sgdma_mm2s_m_read_read                                : in  std_logic                     := 'X';             -- read
			sgdma_mm2s_m_read_readdata                            : out std_logic_vector(7 downto 0);                     -- readdata
			sgdma_mm2s_m_read_readdatavalid                       : out std_logic;                                        -- readdatavalid
			sgdma_s2mm_descriptor_read_address                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_s2mm_descriptor_read_waitrequest                : out std_logic;                                        -- waitrequest
			sgdma_s2mm_descriptor_read_read                       : in  std_logic                     := 'X';             -- read
			sgdma_s2mm_descriptor_read_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			sgdma_s2mm_descriptor_read_readdatavalid              : out std_logic;                                        -- readdatavalid
			sgdma_s2mm_descriptor_write_address                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_s2mm_descriptor_write_waitrequest               : out std_logic;                                        -- waitrequest
			sgdma_s2mm_descriptor_write_write                     : in  std_logic                     := 'X';             -- write
			sgdma_s2mm_descriptor_write_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sgdma_s2mm_m_write_address                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_s2mm_m_write_waitrequest                        : out std_logic;                                        -- waitrequest
			sgdma_s2mm_m_write_byteenable                         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			sgdma_s2mm_m_write_write                              : in  std_logic                     := 'X';             -- write
			sgdma_s2mm_m_write_writedata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			histeq_calc_0_params_address                          : out std_logic_vector(0 downto 0);                     -- address
			histeq_calc_0_params_write                            : out std_logic;                                        -- write
			histeq_calc_0_params_read                             : out std_logic;                                        -- read
			histeq_calc_0_params_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			histeq_calc_0_params_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			histeq_calc_0_params_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_address                 : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                   : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                    : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest             : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect              : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                  : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                    : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                     : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable               : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest              : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess              : out std_logic;                                        -- debugaccess
			performance_counter_0_control_slave_address           : out std_logic_vector(3 downto 0);                     -- address
			performance_counter_0_control_slave_write             : out std_logic;                                        -- write
			performance_counter_0_control_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			performance_counter_0_control_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			performance_counter_0_control_slave_begintransfer     : out std_logic;                                        -- begintransfer
			pll_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pll_pll_slave_write                                   : out std_logic;                                        -- write
			pll_pll_slave_read                                    : out std_logic;                                        -- read
			pll_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_s1_address                                      : out std_logic_vector(23 downto 0);                    -- address
			sdram_s1_write                                        : out std_logic;                                        -- write
			sdram_s1_read                                         : out std_logic;                                        -- read
			sdram_s1_readdata                                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                                    : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                                   : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                                   : out std_logic;                                        -- chipselect
			sgdma_mm2s_csr_address                                : out std_logic_vector(3 downto 0);                     -- address
			sgdma_mm2s_csr_write                                  : out std_logic;                                        -- write
			sgdma_mm2s_csr_read                                   : out std_logic;                                        -- read
			sgdma_mm2s_csr_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sgdma_mm2s_csr_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			sgdma_mm2s_csr_chipselect                             : out std_logic;                                        -- chipselect
			sgdma_s2mm_csr_address                                : out std_logic_vector(3 downto 0);                     -- address
			sgdma_s2mm_csr_write                                  : out std_logic;                                        -- write
			sgdma_s2mm_csr_read                                   : out std_logic;                                        -- read
			sgdma_s2mm_csr_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sgdma_s2mm_csr_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			sgdma_s2mm_csr_chipselect                             : out std_logic                                         -- chipselect
		);
	end component processor_system_mm_interconnect_0;

	component processor_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component processor_system_irq_mapper;

	component processor_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component processor_system_rst_controller;

	component processor_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component processor_system_rst_controller_001;

	signal sgdma_mm2s_out_valid                                                : std_logic;                     -- sgdma_mm2s:out_valid -> histeq_calc_0:asi_in_valid
	signal sgdma_mm2s_out_data                                                 : std_logic_vector(7 downto 0);  -- sgdma_mm2s:out_data -> histeq_calc_0:asi_in_data
	signal sgdma_mm2s_out_ready                                                : std_logic;                     -- histeq_calc_0:asi_in_ready -> sgdma_mm2s:out_ready
	signal sgdma_mm2s_out_startofpacket                                        : std_logic;                     -- sgdma_mm2s:out_startofpacket -> histeq_calc_0:asi_in_sop
	signal sgdma_mm2s_out_endofpacket                                          : std_logic;                     -- sgdma_mm2s:out_endofpacket -> histeq_calc_0:asi_in_eop
	signal histeq_calc_0_out_valid                                             : std_logic;                     -- histeq_calc_0:aso_out_valid -> sgdma_s2mm:in_valid
	signal histeq_calc_0_out_data                                              : std_logic_vector(31 downto 0); -- histeq_calc_0:aso_out_data -> sgdma_s2mm:in_data
	signal histeq_calc_0_out_ready                                             : std_logic;                     -- sgdma_s2mm:in_ready -> histeq_calc_0:aso_out_ready
	signal histeq_calc_0_out_startofpacket                                     : std_logic;                     -- histeq_calc_0:aso_out_sop -> sgdma_s2mm:in_startofpacket
	signal histeq_calc_0_out_endofpacket                                       : std_logic;                     -- histeq_calc_0:aso_out_eop -> sgdma_s2mm:in_endofpacket
	signal histeq_calc_0_out_empty                                             : std_logic;                     -- histeq_calc_0:aso_out_empty -> sgdma_s2mm:in_empty
	signal pll_c0_clk                                                          : std_logic;                     -- pll:c0 -> [histeq_calc_0:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:pll_c0_clk, nios2_gen2_0:clk, performance_counter_0:clk, rst_controller:clk, sdram:clk, sgdma_mm2s:clk, sgdma_s2mm:clk]
	signal nios2_gen2_0_data_master_readdata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                    : std_logic_vector(26 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                 : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                       : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                      : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                  : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal sgdma_mm2s_descriptor_read_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_mm2s_descriptor_read_readdata -> sgdma_mm2s:descriptor_read_readdata
	signal sgdma_mm2s_descriptor_read_waitrequest                              : std_logic;                     -- mm_interconnect_0:sgdma_mm2s_descriptor_read_waitrequest -> sgdma_mm2s:descriptor_read_waitrequest
	signal sgdma_mm2s_descriptor_read_address                                  : std_logic_vector(31 downto 0); -- sgdma_mm2s:descriptor_read_address -> mm_interconnect_0:sgdma_mm2s_descriptor_read_address
	signal sgdma_mm2s_descriptor_read_read                                     : std_logic;                     -- sgdma_mm2s:descriptor_read_read -> mm_interconnect_0:sgdma_mm2s_descriptor_read_read
	signal sgdma_mm2s_descriptor_read_readdatavalid                            : std_logic;                     -- mm_interconnect_0:sgdma_mm2s_descriptor_read_readdatavalid -> sgdma_mm2s:descriptor_read_readdatavalid
	signal sgdma_s2mm_descriptor_read_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_s2mm_descriptor_read_readdata -> sgdma_s2mm:descriptor_read_readdata
	signal sgdma_s2mm_descriptor_read_waitrequest                              : std_logic;                     -- mm_interconnect_0:sgdma_s2mm_descriptor_read_waitrequest -> sgdma_s2mm:descriptor_read_waitrequest
	signal sgdma_s2mm_descriptor_read_address                                  : std_logic_vector(31 downto 0); -- sgdma_s2mm:descriptor_read_address -> mm_interconnect_0:sgdma_s2mm_descriptor_read_address
	signal sgdma_s2mm_descriptor_read_read                                     : std_logic;                     -- sgdma_s2mm:descriptor_read_read -> mm_interconnect_0:sgdma_s2mm_descriptor_read_read
	signal sgdma_s2mm_descriptor_read_readdatavalid                            : std_logic;                     -- mm_interconnect_0:sgdma_s2mm_descriptor_read_readdatavalid -> sgdma_s2mm:descriptor_read_readdatavalid
	signal sgdma_mm2s_descriptor_write_waitrequest                             : std_logic;                     -- mm_interconnect_0:sgdma_mm2s_descriptor_write_waitrequest -> sgdma_mm2s:descriptor_write_waitrequest
	signal sgdma_mm2s_descriptor_write_address                                 : std_logic_vector(31 downto 0); -- sgdma_mm2s:descriptor_write_address -> mm_interconnect_0:sgdma_mm2s_descriptor_write_address
	signal sgdma_mm2s_descriptor_write_write                                   : std_logic;                     -- sgdma_mm2s:descriptor_write_write -> mm_interconnect_0:sgdma_mm2s_descriptor_write_write
	signal sgdma_mm2s_descriptor_write_writedata                               : std_logic_vector(31 downto 0); -- sgdma_mm2s:descriptor_write_writedata -> mm_interconnect_0:sgdma_mm2s_descriptor_write_writedata
	signal sgdma_s2mm_descriptor_write_waitrequest                             : std_logic;                     -- mm_interconnect_0:sgdma_s2mm_descriptor_write_waitrequest -> sgdma_s2mm:descriptor_write_waitrequest
	signal sgdma_s2mm_descriptor_write_address                                 : std_logic_vector(31 downto 0); -- sgdma_s2mm:descriptor_write_address -> mm_interconnect_0:sgdma_s2mm_descriptor_write_address
	signal sgdma_s2mm_descriptor_write_write                                   : std_logic;                     -- sgdma_s2mm:descriptor_write_write -> mm_interconnect_0:sgdma_s2mm_descriptor_write_write
	signal sgdma_s2mm_descriptor_write_writedata                               : std_logic_vector(31 downto 0); -- sgdma_s2mm:descriptor_write_writedata -> mm_interconnect_0:sgdma_s2mm_descriptor_write_writedata
	signal nios2_gen2_0_instruction_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                             : std_logic_vector(26 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal sgdma_mm2s_m_read_readdata                                          : std_logic_vector(7 downto 0);  -- mm_interconnect_0:sgdma_mm2s_m_read_readdata -> sgdma_mm2s:m_read_readdata
	signal sgdma_mm2s_m_read_waitrequest                                       : std_logic;                     -- mm_interconnect_0:sgdma_mm2s_m_read_waitrequest -> sgdma_mm2s:m_read_waitrequest
	signal sgdma_mm2s_m_read_address                                           : std_logic_vector(31 downto 0); -- sgdma_mm2s:m_read_address -> mm_interconnect_0:sgdma_mm2s_m_read_address
	signal sgdma_mm2s_m_read_read                                              : std_logic;                     -- sgdma_mm2s:m_read_read -> mm_interconnect_0:sgdma_mm2s_m_read_read
	signal sgdma_mm2s_m_read_readdatavalid                                     : std_logic;                     -- mm_interconnect_0:sgdma_mm2s_m_read_readdatavalid -> sgdma_mm2s:m_read_readdatavalid
	signal sgdma_s2mm_m_write_waitrequest                                      : std_logic;                     -- mm_interconnect_0:sgdma_s2mm_m_write_waitrequest -> sgdma_s2mm:m_write_waitrequest
	signal sgdma_s2mm_m_write_address                                          : std_logic_vector(31 downto 0); -- sgdma_s2mm:m_write_address -> mm_interconnect_0:sgdma_s2mm_m_write_address
	signal sgdma_s2mm_m_write_byteenable                                       : std_logic_vector(3 downto 0);  -- sgdma_s2mm:m_write_byteenable -> mm_interconnect_0:sgdma_s2mm_m_write_byteenable
	signal sgdma_s2mm_m_write_write                                            : std_logic;                     -- sgdma_s2mm:m_write_write -> mm_interconnect_0:sgdma_s2mm_m_write_write
	signal sgdma_s2mm_m_write_writedata                                        : std_logic_vector(31 downto 0); -- sgdma_s2mm:m_write_writedata -> mm_interconnect_0:sgdma_s2mm_m_write_writedata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect          : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata            : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest         : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write               : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_performance_counter_0_control_slave_readdata      : std_logic_vector(31 downto 0); -- performance_counter_0:readdata -> mm_interconnect_0:performance_counter_0_control_slave_readdata
	signal mm_interconnect_0_performance_counter_0_control_slave_address       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:performance_counter_0_control_slave_address -> performance_counter_0:address
	signal mm_interconnect_0_performance_counter_0_control_slave_begintransfer : std_logic;                     -- mm_interconnect_0:performance_counter_0_control_slave_begintransfer -> performance_counter_0:begintransfer
	signal mm_interconnect_0_performance_counter_0_control_slave_write         : std_logic;                     -- mm_interconnect_0:performance_counter_0_control_slave_write -> performance_counter_0:write
	signal mm_interconnect_0_performance_counter_0_control_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:performance_counter_0_control_slave_writedata -> performance_counter_0:writedata
	signal mm_interconnect_0_sgdma_mm2s_csr_chipselect                         : std_logic;                     -- mm_interconnect_0:sgdma_mm2s_csr_chipselect -> sgdma_mm2s:csr_chipselect
	signal mm_interconnect_0_sgdma_mm2s_csr_readdata                           : std_logic_vector(31 downto 0); -- sgdma_mm2s:csr_readdata -> mm_interconnect_0:sgdma_mm2s_csr_readdata
	signal mm_interconnect_0_sgdma_mm2s_csr_address                            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sgdma_mm2s_csr_address -> sgdma_mm2s:csr_address
	signal mm_interconnect_0_sgdma_mm2s_csr_read                               : std_logic;                     -- mm_interconnect_0:sgdma_mm2s_csr_read -> sgdma_mm2s:csr_read
	signal mm_interconnect_0_sgdma_mm2s_csr_write                              : std_logic;                     -- mm_interconnect_0:sgdma_mm2s_csr_write -> sgdma_mm2s:csr_write
	signal mm_interconnect_0_sgdma_mm2s_csr_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_mm2s_csr_writedata -> sgdma_mm2s:csr_writedata
	signal mm_interconnect_0_sgdma_s2mm_csr_chipselect                         : std_logic;                     -- mm_interconnect_0:sgdma_s2mm_csr_chipselect -> sgdma_s2mm:csr_chipselect
	signal mm_interconnect_0_sgdma_s2mm_csr_readdata                           : std_logic_vector(31 downto 0); -- sgdma_s2mm:csr_readdata -> mm_interconnect_0:sgdma_s2mm_csr_readdata
	signal mm_interconnect_0_sgdma_s2mm_csr_address                            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sgdma_s2mm_csr_address -> sgdma_s2mm:csr_address
	signal mm_interconnect_0_sgdma_s2mm_csr_read                               : std_logic;                     -- mm_interconnect_0:sgdma_s2mm_csr_read -> sgdma_s2mm:csr_read
	signal mm_interconnect_0_sgdma_s2mm_csr_write                              : std_logic;                     -- mm_interconnect_0:sgdma_s2mm_csr_write -> sgdma_s2mm:csr_write
	signal mm_interconnect_0_sgdma_s2mm_csr_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_s2mm_csr_writedata -> sgdma_s2mm:csr_writedata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata             : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest          : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess          : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address              : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read                 : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write                : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_histeq_calc_0_params_readdata                     : std_logic_vector(31 downto 0); -- histeq_calc_0:avs_params_readdata -> mm_interconnect_0:histeq_calc_0_params_readdata
	signal mm_interconnect_0_histeq_calc_0_params_waitrequest                  : std_logic;                     -- histeq_calc_0:avs_params_waitrequest -> mm_interconnect_0:histeq_calc_0_params_waitrequest
	signal mm_interconnect_0_histeq_calc_0_params_address                      : std_logic_vector(0 downto 0);  -- mm_interconnect_0:histeq_calc_0_params_address -> histeq_calc_0:avs_params_address
	signal mm_interconnect_0_histeq_calc_0_params_read                         : std_logic;                     -- mm_interconnect_0:histeq_calc_0_params_read -> histeq_calc_0:avs_params_read
	signal mm_interconnect_0_histeq_calc_0_params_write                        : std_logic;                     -- mm_interconnect_0:histeq_calc_0_params_write -> histeq_calc_0:avs_params_write
	signal mm_interconnect_0_histeq_calc_0_params_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:histeq_calc_0_params_writedata -> histeq_calc_0:avs_params_writedata
	signal mm_interconnect_0_pll_pll_slave_readdata                            : std_logic_vector(31 downto 0); -- pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	signal mm_interconnect_0_pll_pll_slave_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pll_pll_slave_address -> pll:address
	signal mm_interconnect_0_pll_pll_slave_read                                : std_logic;                     -- mm_interconnect_0:pll_pll_slave_read -> pll:read
	signal mm_interconnect_0_pll_pll_slave_write                               : std_logic;                     -- mm_interconnect_0:pll_pll_slave_write -> pll:write
	signal mm_interconnect_0_pll_pll_slave_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	signal mm_interconnect_0_sdram_s1_chipselect                               : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                                 : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                              : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                                  : std_logic_vector(23 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                                     : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                            : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                    : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                                : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal irq_mapper_receiver0_irq                                            : std_logic;                     -- sgdma_mm2s:csr_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                            : std_logic;                     -- sgdma_s2mm:csr_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                            : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver2_irq
	signal nios2_gen2_0_irq_irq                                                : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                      : std_logic;                     -- rst_controller:reset_out -> [histeq_calc_0:reset, irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                  : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	signal nios2_gen2_0_debug_reset_request_reset                              : std_logic;                     -- nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                                  : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]
	signal reset_reset_n_ports_inv                                             : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv      : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv     : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                           : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                          : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                            : std_logic;                     -- rst_controller_reset_out_reset:inv -> [jtag_uart_0:rst_n, nios2_gen2_0:reset_n, performance_counter_0:reset_n, sdram:reset_n, sgdma_mm2s:system_reset_n, sgdma_s2mm:system_reset_n]

begin

	histeq_calc_0 : component acc_linear_function
		port map (
			reset                  => rst_controller_reset_out_reset,                     --  reset.reset
			avs_params_address     => mm_interconnect_0_histeq_calc_0_params_address(0),  -- params.address
			avs_params_read        => mm_interconnect_0_histeq_calc_0_params_read,        --       .read
			avs_params_readdata    => mm_interconnect_0_histeq_calc_0_params_readdata,    --       .readdata
			avs_params_write       => mm_interconnect_0_histeq_calc_0_params_write,       --       .write
			avs_params_writedata   => mm_interconnect_0_histeq_calc_0_params_writedata,   --       .writedata
			avs_params_waitrequest => mm_interconnect_0_histeq_calc_0_params_waitrequest, --       .waitrequest
			clk                    => pll_c0_clk,                                         --  clock.clk
			asi_in_data            => sgdma_mm2s_out_data,                                --     in.data
			asi_in_ready           => sgdma_mm2s_out_ready,                               --       .ready
			asi_in_valid           => sgdma_mm2s_out_valid,                               --       .valid
			asi_in_eop             => sgdma_mm2s_out_endofpacket,                         --       .endofpacket
			asi_in_sop             => sgdma_mm2s_out_startofpacket,                       --       .startofpacket
			aso_out_data           => histeq_calc_0_out_data,                             --    out.data
			aso_out_ready          => histeq_calc_0_out_ready,                            --       .ready
			aso_out_valid          => histeq_calc_0_out_valid,                            --       .valid
			aso_out_empty          => histeq_calc_0_out_empty,                            --       .empty
			aso_out_eop            => histeq_calc_0_out_endofpacket,                      --       .endofpacket
			aso_out_sop            => histeq_calc_0_out_startofpacket                     --       .startofpacket
		);

	jtag_uart_0 : component processor_system_jtag_uart_0
		port map (
			clk            => pll_c0_clk,                                                      --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver2_irq                                         --               irq.irq
		);

	nios2_gen2_0 : component processor_system_nios2_gen2_0
		port map (
			clk                                 => pll_c0_clk,                                                 --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	performance_counter_0 : component processor_system_performance_counter_0
		port map (
			clk           => pll_c0_clk,                                                          --           clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                            --         reset.reset_n
			address       => mm_interconnect_0_performance_counter_0_control_slave_address,       -- control_slave.address
			begintransfer => mm_interconnect_0_performance_counter_0_control_slave_begintransfer, --              .begintransfer
			readdata      => mm_interconnect_0_performance_counter_0_control_slave_readdata,      --              .readdata
			write         => mm_interconnect_0_performance_counter_0_control_slave_write,         --              .write
			writedata     => mm_interconnect_0_performance_counter_0_control_slave_writedata      --              .writedata
		);

	pll : component processor_system_pll
		port map (
			clk                => clk_clk,                                   --       inclk_interface.clk
			reset              => rst_controller_001_reset_out_reset,        -- inclk_interface_reset.reset
			read               => mm_interconnect_0_pll_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_pll_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_pll_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_pll_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_pll_pll_slave_writedata, --                      .writedata
			c0                 => pll_c0_clk,                                --                    c0.clk
			c1                 => sdram_clk_clk,                             --                    c1.clk
			scandone           => open,                                      --           (terminated)
			scandataout        => open,                                      --           (terminated)
			areset             => '0',                                       --           (terminated)
			locked             => open,                                      --           (terminated)
			phasedone          => open,                                      --           (terminated)
			phasecounterselect => "0000",                                    --           (terminated)
			phaseupdown        => '0',                                       --           (terminated)
			phasestep          => '0',                                       --           (terminated)
			scanclk            => '0',                                       --           (terminated)
			scanclkena         => '0',                                       --           (terminated)
			scandata           => '0',                                       --           (terminated)
			configupdate       => '0'                                        --           (terminated)
		);

	sdram : component processor_system_sdram
		port map (
			clk            => pll_c0_clk,                                      --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	sgdma_mm2s : component processor_system_sgdma_mm2s
		port map (
			clk                           => pll_c0_clk,                                  --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv,    --            reset.reset_n
			csr_chipselect                => mm_interconnect_0_sgdma_mm2s_csr_chipselect, --              csr.chipselect
			csr_address                   => mm_interconnect_0_sgdma_mm2s_csr_address,    --                 .address
			csr_read                      => mm_interconnect_0_sgdma_mm2s_csr_read,       --                 .read
			csr_write                     => mm_interconnect_0_sgdma_mm2s_csr_write,      --                 .write
			csr_writedata                 => mm_interconnect_0_sgdma_mm2s_csr_writedata,  --                 .writedata
			csr_readdata                  => mm_interconnect_0_sgdma_mm2s_csr_readdata,   --                 .readdata
			descriptor_read_readdata      => sgdma_mm2s_descriptor_read_readdata,         --  descriptor_read.readdata
			descriptor_read_readdatavalid => sgdma_mm2s_descriptor_read_readdatavalid,    --                 .readdatavalid
			descriptor_read_waitrequest   => sgdma_mm2s_descriptor_read_waitrequest,      --                 .waitrequest
			descriptor_read_address       => sgdma_mm2s_descriptor_read_address,          --                 .address
			descriptor_read_read          => sgdma_mm2s_descriptor_read_read,             --                 .read
			descriptor_write_waitrequest  => sgdma_mm2s_descriptor_write_waitrequest,     -- descriptor_write.waitrequest
			descriptor_write_address      => sgdma_mm2s_descriptor_write_address,         --                 .address
			descriptor_write_write        => sgdma_mm2s_descriptor_write_write,           --                 .write
			descriptor_write_writedata    => sgdma_mm2s_descriptor_write_writedata,       --                 .writedata
			csr_irq                       => irq_mapper_receiver0_irq,                    --          csr_irq.irq
			m_read_readdata               => sgdma_mm2s_m_read_readdata,                  --           m_read.readdata
			m_read_readdatavalid          => sgdma_mm2s_m_read_readdatavalid,             --                 .readdatavalid
			m_read_waitrequest            => sgdma_mm2s_m_read_waitrequest,               --                 .waitrequest
			m_read_address                => sgdma_mm2s_m_read_address,                   --                 .address
			m_read_read                   => sgdma_mm2s_m_read_read,                      --                 .read
			out_data                      => sgdma_mm2s_out_data,                         --              out.data
			out_valid                     => sgdma_mm2s_out_valid,                        --                 .valid
			out_ready                     => sgdma_mm2s_out_ready,                        --                 .ready
			out_endofpacket               => sgdma_mm2s_out_endofpacket,                  --                 .endofpacket
			out_startofpacket             => sgdma_mm2s_out_startofpacket                 --                 .startofpacket
		);

	sgdma_s2mm : component processor_system_sgdma_s2mm
		port map (
			clk                           => pll_c0_clk,                                  --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv,    --            reset.reset_n
			csr_chipselect                => mm_interconnect_0_sgdma_s2mm_csr_chipselect, --              csr.chipselect
			csr_address                   => mm_interconnect_0_sgdma_s2mm_csr_address,    --                 .address
			csr_read                      => mm_interconnect_0_sgdma_s2mm_csr_read,       --                 .read
			csr_write                     => mm_interconnect_0_sgdma_s2mm_csr_write,      --                 .write
			csr_writedata                 => mm_interconnect_0_sgdma_s2mm_csr_writedata,  --                 .writedata
			csr_readdata                  => mm_interconnect_0_sgdma_s2mm_csr_readdata,   --                 .readdata
			descriptor_read_readdata      => sgdma_s2mm_descriptor_read_readdata,         --  descriptor_read.readdata
			descriptor_read_readdatavalid => sgdma_s2mm_descriptor_read_readdatavalid,    --                 .readdatavalid
			descriptor_read_waitrequest   => sgdma_s2mm_descriptor_read_waitrequest,      --                 .waitrequest
			descriptor_read_address       => sgdma_s2mm_descriptor_read_address,          --                 .address
			descriptor_read_read          => sgdma_s2mm_descriptor_read_read,             --                 .read
			descriptor_write_waitrequest  => sgdma_s2mm_descriptor_write_waitrequest,     -- descriptor_write.waitrequest
			descriptor_write_address      => sgdma_s2mm_descriptor_write_address,         --                 .address
			descriptor_write_write        => sgdma_s2mm_descriptor_write_write,           --                 .write
			descriptor_write_writedata    => sgdma_s2mm_descriptor_write_writedata,       --                 .writedata
			csr_irq                       => irq_mapper_receiver1_irq,                    --          csr_irq.irq
			in_startofpacket              => histeq_calc_0_out_startofpacket,             --               in.startofpacket
			in_endofpacket                => histeq_calc_0_out_endofpacket,               --                 .endofpacket
			in_data                       => histeq_calc_0_out_data,                      --                 .data
			in_valid                      => histeq_calc_0_out_valid,                     --                 .valid
			in_ready                      => histeq_calc_0_out_ready,                     --                 .ready
			in_empty                      => histeq_calc_0_out_empty,                     --                 .empty
			m_write_waitrequest           => sgdma_s2mm_m_write_waitrequest,              --          m_write.waitrequest
			m_write_address               => sgdma_s2mm_m_write_address,                  --                 .address
			m_write_write                 => sgdma_s2mm_m_write_write,                    --                 .write
			m_write_writedata             => sgdma_s2mm_m_write_writedata,                --                 .writedata
			m_write_byteenable            => sgdma_s2mm_m_write_byteenable                --                 .byteenable
		);

	mm_interconnect_0 : component processor_system_mm_interconnect_0
		port map (
			clk_0_clk_clk                                         => clk_clk,                                                             --                                       clk_0_clk.clk
			pll_c0_clk                                            => pll_c0_clk,                                                          --                                          pll_c0.clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset        => rst_controller_reset_out_reset,                                      --        nios2_gen2_0_reset_reset_bridge_in_reset.reset
			pll_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                                  -- pll_inclk_interface_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                      => nios2_gen2_0_data_master_address,                                    --                        nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                  => nios2_gen2_0_data_master_waitrequest,                                --                                                .waitrequest
			nios2_gen2_0_data_master_byteenable                   => nios2_gen2_0_data_master_byteenable,                                 --                                                .byteenable
			nios2_gen2_0_data_master_read                         => nios2_gen2_0_data_master_read,                                       --                                                .read
			nios2_gen2_0_data_master_readdata                     => nios2_gen2_0_data_master_readdata,                                   --                                                .readdata
			nios2_gen2_0_data_master_write                        => nios2_gen2_0_data_master_write,                                      --                                                .write
			nios2_gen2_0_data_master_writedata                    => nios2_gen2_0_data_master_writedata,                                  --                                                .writedata
			nios2_gen2_0_data_master_debugaccess                  => nios2_gen2_0_data_master_debugaccess,                                --                                                .debugaccess
			nios2_gen2_0_instruction_master_address               => nios2_gen2_0_instruction_master_address,                             --                 nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest           => nios2_gen2_0_instruction_master_waitrequest,                         --                                                .waitrequest
			nios2_gen2_0_instruction_master_read                  => nios2_gen2_0_instruction_master_read,                                --                                                .read
			nios2_gen2_0_instruction_master_readdata              => nios2_gen2_0_instruction_master_readdata,                            --                                                .readdata
			sgdma_mm2s_descriptor_read_address                    => sgdma_mm2s_descriptor_read_address,                                  --                      sgdma_mm2s_descriptor_read.address
			sgdma_mm2s_descriptor_read_waitrequest                => sgdma_mm2s_descriptor_read_waitrequest,                              --                                                .waitrequest
			sgdma_mm2s_descriptor_read_read                       => sgdma_mm2s_descriptor_read_read,                                     --                                                .read
			sgdma_mm2s_descriptor_read_readdata                   => sgdma_mm2s_descriptor_read_readdata,                                 --                                                .readdata
			sgdma_mm2s_descriptor_read_readdatavalid              => sgdma_mm2s_descriptor_read_readdatavalid,                            --                                                .readdatavalid
			sgdma_mm2s_descriptor_write_address                   => sgdma_mm2s_descriptor_write_address,                                 --                     sgdma_mm2s_descriptor_write.address
			sgdma_mm2s_descriptor_write_waitrequest               => sgdma_mm2s_descriptor_write_waitrequest,                             --                                                .waitrequest
			sgdma_mm2s_descriptor_write_write                     => sgdma_mm2s_descriptor_write_write,                                   --                                                .write
			sgdma_mm2s_descriptor_write_writedata                 => sgdma_mm2s_descriptor_write_writedata,                               --                                                .writedata
			sgdma_mm2s_m_read_address                             => sgdma_mm2s_m_read_address,                                           --                               sgdma_mm2s_m_read.address
			sgdma_mm2s_m_read_waitrequest                         => sgdma_mm2s_m_read_waitrequest,                                       --                                                .waitrequest
			sgdma_mm2s_m_read_read                                => sgdma_mm2s_m_read_read,                                              --                                                .read
			sgdma_mm2s_m_read_readdata                            => sgdma_mm2s_m_read_readdata,                                          --                                                .readdata
			sgdma_mm2s_m_read_readdatavalid                       => sgdma_mm2s_m_read_readdatavalid,                                     --                                                .readdatavalid
			sgdma_s2mm_descriptor_read_address                    => sgdma_s2mm_descriptor_read_address,                                  --                      sgdma_s2mm_descriptor_read.address
			sgdma_s2mm_descriptor_read_waitrequest                => sgdma_s2mm_descriptor_read_waitrequest,                              --                                                .waitrequest
			sgdma_s2mm_descriptor_read_read                       => sgdma_s2mm_descriptor_read_read,                                     --                                                .read
			sgdma_s2mm_descriptor_read_readdata                   => sgdma_s2mm_descriptor_read_readdata,                                 --                                                .readdata
			sgdma_s2mm_descriptor_read_readdatavalid              => sgdma_s2mm_descriptor_read_readdatavalid,                            --                                                .readdatavalid
			sgdma_s2mm_descriptor_write_address                   => sgdma_s2mm_descriptor_write_address,                                 --                     sgdma_s2mm_descriptor_write.address
			sgdma_s2mm_descriptor_write_waitrequest               => sgdma_s2mm_descriptor_write_waitrequest,                             --                                                .waitrequest
			sgdma_s2mm_descriptor_write_write                     => sgdma_s2mm_descriptor_write_write,                                   --                                                .write
			sgdma_s2mm_descriptor_write_writedata                 => sgdma_s2mm_descriptor_write_writedata,                               --                                                .writedata
			sgdma_s2mm_m_write_address                            => sgdma_s2mm_m_write_address,                                          --                              sgdma_s2mm_m_write.address
			sgdma_s2mm_m_write_waitrequest                        => sgdma_s2mm_m_write_waitrequest,                                      --                                                .waitrequest
			sgdma_s2mm_m_write_byteenable                         => sgdma_s2mm_m_write_byteenable,                                       --                                                .byteenable
			sgdma_s2mm_m_write_write                              => sgdma_s2mm_m_write_write,                                            --                                                .write
			sgdma_s2mm_m_write_writedata                          => sgdma_s2mm_m_write_writedata,                                        --                                                .writedata
			histeq_calc_0_params_address                          => mm_interconnect_0_histeq_calc_0_params_address,                      --                            histeq_calc_0_params.address
			histeq_calc_0_params_write                            => mm_interconnect_0_histeq_calc_0_params_write,                        --                                                .write
			histeq_calc_0_params_read                             => mm_interconnect_0_histeq_calc_0_params_read,                         --                                                .read
			histeq_calc_0_params_readdata                         => mm_interconnect_0_histeq_calc_0_params_readdata,                     --                                                .readdata
			histeq_calc_0_params_writedata                        => mm_interconnect_0_histeq_calc_0_params_writedata,                    --                                                .writedata
			histeq_calc_0_params_waitrequest                      => mm_interconnect_0_histeq_calc_0_params_waitrequest,                  --                                                .waitrequest
			jtag_uart_0_avalon_jtag_slave_address                 => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,             --                   jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,               --                                                .write
			jtag_uart_0_avalon_jtag_slave_read                    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,                --                                                .read
			jtag_uart_0_avalon_jtag_slave_readdata                => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,            --                                                .readdata
			jtag_uart_0_avalon_jtag_slave_writedata               => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,           --                                                .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,         --                                                .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect              => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,          --                                                .chipselect
			nios2_gen2_0_debug_mem_slave_address                  => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,              --                    nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                    => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,                --                                                .write
			nios2_gen2_0_debug_mem_slave_read                     => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,                 --                                                .read
			nios2_gen2_0_debug_mem_slave_readdata                 => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,             --                                                .readdata
			nios2_gen2_0_debug_mem_slave_writedata                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,            --                                                .writedata
			nios2_gen2_0_debug_mem_slave_byteenable               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,           --                                                .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,          --                                                .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,          --                                                .debugaccess
			performance_counter_0_control_slave_address           => mm_interconnect_0_performance_counter_0_control_slave_address,       --             performance_counter_0_control_slave.address
			performance_counter_0_control_slave_write             => mm_interconnect_0_performance_counter_0_control_slave_write,         --                                                .write
			performance_counter_0_control_slave_readdata          => mm_interconnect_0_performance_counter_0_control_slave_readdata,      --                                                .readdata
			performance_counter_0_control_slave_writedata         => mm_interconnect_0_performance_counter_0_control_slave_writedata,     --                                                .writedata
			performance_counter_0_control_slave_begintransfer     => mm_interconnect_0_performance_counter_0_control_slave_begintransfer, --                                                .begintransfer
			pll_pll_slave_address                                 => mm_interconnect_0_pll_pll_slave_address,                             --                                   pll_pll_slave.address
			pll_pll_slave_write                                   => mm_interconnect_0_pll_pll_slave_write,                               --                                                .write
			pll_pll_slave_read                                    => mm_interconnect_0_pll_pll_slave_read,                                --                                                .read
			pll_pll_slave_readdata                                => mm_interconnect_0_pll_pll_slave_readdata,                            --                                                .readdata
			pll_pll_slave_writedata                               => mm_interconnect_0_pll_pll_slave_writedata,                           --                                                .writedata
			sdram_s1_address                                      => mm_interconnect_0_sdram_s1_address,                                  --                                        sdram_s1.address
			sdram_s1_write                                        => mm_interconnect_0_sdram_s1_write,                                    --                                                .write
			sdram_s1_read                                         => mm_interconnect_0_sdram_s1_read,                                     --                                                .read
			sdram_s1_readdata                                     => mm_interconnect_0_sdram_s1_readdata,                                 --                                                .readdata
			sdram_s1_writedata                                    => mm_interconnect_0_sdram_s1_writedata,                                --                                                .writedata
			sdram_s1_byteenable                                   => mm_interconnect_0_sdram_s1_byteenable,                               --                                                .byteenable
			sdram_s1_readdatavalid                                => mm_interconnect_0_sdram_s1_readdatavalid,                            --                                                .readdatavalid
			sdram_s1_waitrequest                                  => mm_interconnect_0_sdram_s1_waitrequest,                              --                                                .waitrequest
			sdram_s1_chipselect                                   => mm_interconnect_0_sdram_s1_chipselect,                               --                                                .chipselect
			sgdma_mm2s_csr_address                                => mm_interconnect_0_sgdma_mm2s_csr_address,                            --                                  sgdma_mm2s_csr.address
			sgdma_mm2s_csr_write                                  => mm_interconnect_0_sgdma_mm2s_csr_write,                              --                                                .write
			sgdma_mm2s_csr_read                                   => mm_interconnect_0_sgdma_mm2s_csr_read,                               --                                                .read
			sgdma_mm2s_csr_readdata                               => mm_interconnect_0_sgdma_mm2s_csr_readdata,                           --                                                .readdata
			sgdma_mm2s_csr_writedata                              => mm_interconnect_0_sgdma_mm2s_csr_writedata,                          --                                                .writedata
			sgdma_mm2s_csr_chipselect                             => mm_interconnect_0_sgdma_mm2s_csr_chipselect,                         --                                                .chipselect
			sgdma_s2mm_csr_address                                => mm_interconnect_0_sgdma_s2mm_csr_address,                            --                                  sgdma_s2mm_csr.address
			sgdma_s2mm_csr_write                                  => mm_interconnect_0_sgdma_s2mm_csr_write,                              --                                                .write
			sgdma_s2mm_csr_read                                   => mm_interconnect_0_sgdma_s2mm_csr_read,                               --                                                .read
			sgdma_s2mm_csr_readdata                               => mm_interconnect_0_sgdma_s2mm_csr_readdata,                           --                                                .readdata
			sgdma_s2mm_csr_writedata                              => mm_interconnect_0_sgdma_s2mm_csr_writedata,                          --                                                .writedata
			sgdma_s2mm_csr_chipselect                             => mm_interconnect_0_sgdma_s2mm_csr_chipselect                          --                                                .chipselect
		);

	irq_mapper : component processor_system_irq_mapper
		port map (
			clk           => pll_c0_clk,                     --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component processor_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => pll_c0_clk,                             --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_001 : component processor_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of processor_system
